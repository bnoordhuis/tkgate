//: version "2.0"
//: property title = "edit1_tut.v"
//: property useExtBars = 0
//: property discardChanges = 1

module main;    //: root_module
wire w7;    //: /sn:0 {0}(682,363)(697,363)(697,375){1}
wire s0;    //: {0}(750,310)(780,310){1}
wire w4;    //: /sn:0 {0}(702,345)(702,375){1}
wire c0;    //: {0}(598,268)(704,268)(704,310){1}
//: {2}(706,312)(729,312){3}
//: {4}(704,314)(704,324){5}
wire c1;    //: {0}(700,396)(700,433){1}
//: {2}(702,435)(725,435){3}
//: {4}(700,437)(700,447){5}
wire s1;    //: /dp:1 {0}(746,433)(781,433){1}
wire a1;    //: {0}(598,427)(638,427){1}
//: {2}(642,427)(650,427){3}
//: {4}(640,429)(640,483)(657,483){5}
wire b1;    //: {0}(598,462)(632,462){1}
//: {2}(634,460)(634,432)(650,432){3}
//: {4}(634,464)(634,488)(657,488){5}
wire w8;    //: /sn:0 {0}(678,486)(693,486)(693,498){1}
wire a0;    //: /dp:1 {0}(598,304)(642,304){1}
//: {2}(646,304)(654,304){3}
//: {4}(644,306)(644,360)(661,360){5}
wire b0;    //: /dp:1 {0}(598,339)(636,339){1}
//: {2}(638,337)(638,309)(654,309){3}
//: {4}(638,341)(638,365)(661,365){5}
wire c2;    //: {0}(783,530)(696,530)(696,519){1}
wire w10;    //: /sn:0 {0}(725,430)(697,430){1}
//: {2}(693,430)(671,430){3}
//: {4}(695,432)(695,447){5}
wire w5;    //: /sn:0 {0}(698,468)(698,498){1}
wire w9;    //: /sn:0 {0}(729,307)(701,307){1}
//: {2}(697,307)(675,307){3}
//: {4}(699,309)(699,324){5}
//: enddecls

  //: joint g8 (c1) @(700, 435) /w:[ 2 1 -1 4 ]
  nand g4 (.I0(w8), .I1(w5), .Z(c2));   //: @(696,509) /sn:0 /R:3 /w:[ 1 1 1 ]
  //: comment g61 /dolink:1 /link:"@T/edwire_tut.v" @(622,100) /sn:0
  //: /line:"�磻����Խ�"
  //: /end
  led g37 (.I(s0));   //: @(787,310) /sn:0 /R:3 /w:[ 1 ] /type:0
  xor g34 (.I0(w10), .I1(c1), .Z(s1));   //: @(736,433) /sn:0 /w:[ 0 3 0 ]
  //: comment g3 /dolink:0 /link:"" @(29,249) /anc:1
  //: /line:"5) �֥ġ���ץ�˥塼�Ρ֥ӥå����פ����򤷤ơ���ܥ󥱡��֥�Υġ����Ф�"
  //: /line:"�Ʋ���������������ȡ�������ɥ������ˡ֥ӥå����פ����ϥܥå������Фޤ���"
  //: /line:"�ܥå����򥯥�å����ơ�1��32�ο��������Ϥ��Ʋ����������줫��磻���"
  //: /line:"����å����ơ������Ƥ���ӥå��������ꤷ�ƤߤƲ�������"
  //: /line:""
  //: /line:"6) �֥ġ���ץ�˥塼�Ρְ�ư����³�פ����򤷡��磻�����֥롦����å�����"
  //: /line:"�ȡ�°���ܥå����������ޤ����ͥå�̾���ͥå�̾��ɽ�����뤫�ɤ������ӥå���"
  //: /line:"�ʤɤ�°��������Ǥ��ޤ����ޥ����α��ܥ���Υ�˥塼�Ǥ�����Ǥ��ޤ���"
  //: /line:""
  //: /line:"7) OR�����Ȥʤɤ���֥롦����å�����ȡ������Ȥ�°���ܥå����������ޤ���"
  //: /line:"������̾��������̾��ɽ�����뤫�ɤ����������Ȥ���ư����뤫�ɤ����ʤɤ�"
  //: /line:"°�����������ޤ����ݡ��Ȥ��ɲá�������Խ��ʤɤ����ޤ���"
  //: /line:""
  //: /line:"8) �����Ȥ�ޥ������ܥ���ǥ���å����ơ��ְ�ư�ԲġפΥե饰�򥻥åȤ���"
  //: /line:"�ߤƲ����������Υե饰�����åȤ��Ƥ���С������Ȥΰ�ư�Ͻ���ޤ���"
  //: /end
  //: comment g2 /dolink:0 /link:"" @(29,38) /anc:1
  //: /line:"1) �ޥ����κ��ܥ���ǥ����Ȥ򥯥�å������ܥ���򲡤����ޤ��̤ξ��˰�ư"
  //: /line:"���ƤߤƲ������������Ȥ˷Ҥ��Ǥ���磻�����˰�ư���ޤ���"
  //: /line:""
  //: /line:"2) �֥ġ���ץ�˥塼�Ρ֥磻������ǡפ����򤷤ơ����å����Υġ����"
  //: /line:"�Ф����磻��Τɤ����򥯥�å����ƤߤƲ����������ˤ�Ҥ��Ǥ��ʤ��磻���"
  //: /line:"��ʬ�ϼ�ưŪ�˺������ޤ����ޥ������ܥ���ǳ�����˥塼�����Ѥ��Ƥ�"
  //: /line:"���å�����Ф��ޤ���"
  //: /line:""
  //: /line:"3) �֥ġ���ץ�˥塼�Ρ�����פ����򤷤ơ�����ġ����Ф��������Ȥ�"
  //: /line:"���Ϥ���Ϥ򥯥�å����ƤߤƲ�����������δݤ����줿�ꡢ�ä����ꤷ�ޤ���"
  //: /line:""
  //: /line:"4) �֥ġ���ץ�˥塼�Ρ֥����Ȥκ���פ����򤷡������Ȥ򥯥�å����Ƥߤ�"
  //: /line:"�������������Ȥ��������ޤ��������Ȥ����򤷤ơ��ǥ꡼�ȡ������򲡤����ꡢ"
  //: /line:"�ޥ������ܥ���ǡֺ���פ����򤷤��ꤹ�뤳�ȤǤ⥲���Ȥ�����Ǥ��ޤ���"
  //: /end
  nand g1 (.I0(w7), .I1(w4), .Z(c1));   //: @(700,386) /sn:0 /R:3 /w:[ 1 1 0 ]
  //: switch g11 (a1) @(581,427) /sn:0 /w:[ 0 ] /st:0
  //: comment g16 /dolink:1 /link:"@T/module_tut.v" @(622,115) /sn:0
  //: /line:"�⥸�塼��λȤ���"
  //: /end
  //: joint g10 (a1) @(640, 427) /w:[ 2 -1 1 4 ]
  nand g28 (.I0(a0), .I1(b0), .Z(w7));   //: @(672,363) /sn:0 /w:[ 5 5 0 ]
  led g19 (.I(s1));   //: @(788,433) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: switch g27 (c0) @(581,268) /sn:0 /w:[ 0 ] /st:0
  //: joint g32 (w9) @(699, 307) /w:[ 1 -1 2 4 ]
  //: joint g38 (b1) @(634, 462) /w:[ -1 2 1 4 ]
  nand g6 (.I0(a1), .I1(b1), .Z(w8));   //: @(668,486) /sn:0 /w:[ 5 5 0 ]
  nand g9 (.I0(w10), .I1(c1), .Z(w5));   //: @(698,458) /sn:0 /R:3 /w:[ 5 5 0 ]
  //: joint g7 (w10) @(695, 430) /w:[ 1 -1 2 4 ]
  nand g31 (.I0(w9), .I1(c0), .Z(w4));   //: @(702,335) /sn:0 /R:3 /w:[ 5 5 0 ]
  //: frame g15 @(600,25) /sn:0 /wi:224 /ht:149 /tx:"���塼�ȥꥢ��"
  //: comment g20 /dolink:1 /link:"@T/create_tut.v" @(622,55) /sn:0
  //: /line:"��ϩ�κ���"
  //: /end
  led g39 (.I(c2));   //: @(790,530) /sn:0 /R:3 /w:[ 0 ] /type:0
  //: switch g25 (a0) @(581,304) /sn:0 /w:[ 0 ] /st:0
  //: joint g29 (a0) @(644, 304) /w:[ 2 -1 1 4 ]
  //: comment g17 /dolink:1 /link:"@T/sim_tut.v" @(622,130) /sn:0
  //: /line:"�ȹ礻��ϩ�Υ��ߥ�졼�����"
  //: /end
  //: comment g5 /dolink:0 /link:"@T/edit1_tut.v" @(622,70) /sn:0 /anc:1
  //: /line:"���ܤ��Խ��⡼��"
  //: /end
  //: comment g14 /dolink:1 /link:"@T/seqsim_tut.v" @(622,145) /sn:0
  //: /line:"�����ϩ�Υ��ߥ�졼�����"
  //: /end
  //: switch g36 (b1) @(581,462) /sn:0 /w:[ 0 ] /st:0
  xor g24 (.I0(w9), .I1(c0), .Z(s0));   //: @(740,310) /sn:0 /w:[ 0 3 0 ]
  //: comment g21 /dolink:1 /link:"@T/edit2_tut.v" @(622,85) /sn:0
  //: /line:"���롼�פ��Խ���ǽ"
  //: /end
  xor g23 (.I0(a0), .I1(b0), .Z(w9));   //: @(665,307) /sn:0 /w:[ 3 3 3 ]
  xor g35 (.I0(a1), .I1(b1), .Z(w10));   //: @(661,430) /sn:0 /w:[ 3 3 3 ]
  //: comment g0 /dolink:0 /link:"" @(8,10) /anc:1
  //: /line:"���Υ��塼�ȥꥢ��Ǥϡ�TkGate�δ����Խ���ǽ��Ҳ𤹤롣"
  //: /line:""
  //: /end
  //: switch g26 (b0) @(581,339) /sn:0 /w:[ 0 ] /st:0
  //: comment g22 /dolink:0 /link:"" @(605,70) /sn:0
  //: /line:"->"
  //: /end
  //: comment g18 /dolink:1 /link:"@T/welcome_tut.v" @(622,40) /sn:0
  //: /line:"TkGate�ξҲ�"
  //: /end
  //: joint g30 (b0) @(638, 339) /w:[ -1 2 1 4 ]
  //: joint g33 (c0) @(704, 312) /w:[ 2 1 -1 4 ]

endmodule
