//: version "1.6i"
//: property useExtBars = 0
//: property discardChanges = 1

module main;    //: root_module
wire w32;    //: /sn:0 {0}(631,288)(641,288){1}
wire w6;    //: /sn:0 {0}(484,155)(524,155)(524,138)(549,138)(549,150)(574,150)(574,200)(500,200)(500,170){1}
wire w7;    //: /sn:0 {0}(476,435)(486,435){1}
wire w46;    //: /sn:0 /dp:1 {0}(737,572)(694,572)(694,563){1}
//: {2}(696,561)(710,561)(710,523)(735,523){3}
//: {4}(692,561)(659,561){5}
wire w16;    //: /sn:0 {0}(553,109)(563,109){1}
wire w14;    //: /sn:0 /dp:1 {0}(532,106)(522,106)(522,87)(541,87)(541,54)(488,54){1}
wire w19;    //: /sn:0 {0}(610,437)(620,437){1}
wire w15;    //: /sn:0 {0}(522,111)(532,111){1}
wire w4;    //: /sn:0 {0}(453,157)(463,157){1}
wire w38;    //: /sn:0 {0}(755,394)(765,394){1}
wire w0;    //: /sn:0 {0}(453,152)(463,152){1}
wire w3;    //: /sn:0 {0}(489,288)(530,288){1}
//: {2}(534,288)(587,288){3}
//: {4}(532,286)(532,242)(562,242){5}
wire w37;    //: /sn:0 {0}(729,394)(739,394){1}
wire w34;    //: /sn:0 {0}(752,363)(762,363){1}
wire w43;    //: /sn:0 {0}(628,558)(638,558){1}
wire w21;    //: /sn:0 {0}(610,475)(620,475){1}
wire w31;    //: /sn:0 {0}(631,283)(641,283){1}
wire w28;    //: /sn:0 {0}(662,286)(703,286){1}
//: {2}(707,286)(760,286){3}
//: {4}(705,284)(705,240)(735,240){5}
wire w36;    //: /sn:0 {0}(640,365)(650,365){1}
wire w41;    //: /sn:0 {0}(499,551)(509,551){1}
wire w23;    //: /sn:0 {0}(544,393)(554,393){1}
wire w24;    //: /sn:0 {0}(554,365)(531,365){1}
//: {2}(529,363)(529,334)(555,334){3}
//: {4}(527,365)(489,365){5}
wire w20;    //: /sn:0 {0}(594,475)(582,475)(582,437)(594,437){1}
wire w1;    //: /sn:0 {0}(458,285)(468,285){1}
wire w25;    //: /sn:0 {0}(571,334)(581,334){1}
wire w35;    //: /sn:0 {0}(640,360)(650,360){1}
wire w8;    //: /sn:0 {0}(583,240)(593,240){1}
wire w18;    //: /sn:0 {0}(529,481)(539,481){1}
wire w40;    //: /sn:0 {0}(560,479)(570,479){1}
wire w30;    //: /sn:0 {0}(756,238)(766,238){1}
wire w22;    //: /sn:0 {0}(458,367)(468,367){1}
wire w17;    //: /sn:0 {0}(539,476)(523,476)(523,438)(507,438){1}
wire w44;    //: /sn:0 {0}(628,563)(638,563){1}
wire w12;    //: /sn:0 {0}(457,56)(467,56){1}
wire w11;    //: /sn:0 {0}(457,51)(467,51){1}
wire w2;    //: /sn:0 {0}(458,290)(468,290){1}
wire w10;    //: /sn:0 {0}(458,362)(468,362){1}
wire w13;    //: /sn:0 {0}(499,546)(509,546){1}
wire w27;    //: /sn:0 {0}(570,393)(580,393){1}
wire w48;    //: /sn:0 {0}(751,523)(761,523){1}
wire w33;    //: /sn:0 {0}(736,363)(713,363){1}
//: {2}(711,361)(711,331)(737,331){3}
//: {4}(709,363)(671,363){5}
wire w5;    //: /sn:0 {0}(552,237)(562,237){1}
wire w47;    //: /sn:0 {0}(753,572)(763,572){1}
wire w29;    //: /sn:0 {0}(725,235)(735,235){1}
wire w42;    //: /sn:0 {0}(530,549)(548,549)(548,513){1}
wire w9;    //: /sn:0 {0}(476,440)(486,440){1}
wire w39;    //: /sn:0 {0}(753,331)(763,331){1}
wire w26;    //: /sn:0 {0}(570,365)(580,365){1}
//: enddecls

  //: comment g61 /dolink:0 /link:"@T/edwire_tut.v" @(630,100) /sn:0 /anc:1
  //: /line:"Leitungen editieren"
  //: /end
  xor g8 (.I0(w0), .I1(w4), .Z(w6));   //: @(474,155) /sn:0 /anc:1 /w:[ 1 1 0 ]
  //: comment g4 /dolink:0 /link:"" @(543,256) /sn:0
  //: /line:"<---"
  //: /end
  //: frame g51 @(450,507) /sn:0 /anc:1 /wi:145 /ht:74 /tx:"Bild 6a"
  //: joint g37 (w33) @(711, 363) /w:[ 1 2 4 -1 ]
  //: frame g34 @(449,321) /sn:0 /anc:1 /wi:160 /ht:88 /tx:"Bild 4a"
  //: joint g3 (w3) @(532, 288) /w:[ 2 4 1 -1 ]
  or g13 (.I0(w17), .I1(w18), .Z(w40));   //: @(550,479) /sn:0 /w:[ 0 1 0 ]
  and g2 (.I0(w5), .I1(w3), .Z(w8));   //: @(573,240) /sn:0 /w:[ 1 5 0 ]
  //: comment g1 /dolink:1 /link:"@T/edit1_tut.v" @(630,70) /sn:0 /anc:1
  //: /line:"Grundlegende Editier-Modi"
  //: /end
  and g11 (.I0(w14), .I1(w15), .Z(w16));   //: @(543,109) /sn:0 /anc:1 /w:[ 0 1 0 ]
  //: comment g16 /dolink:1 /link:"@T/module_tut.v" @(630,115) /sn:0 /anc:1
  //: /line:"Module benutzen"
  //: /end
  //: joint g50 (w46) @(694, 561) /w:[ 2 -1 4 1 ]
  buf g28 (.I(w24), .Z(w26));   //: @(560,365) /sn:0 /w:[ 0 0 ]
  and g10 (.I0(w11), .I1(w12), .Z(w14));   //: @(478,54) /sn:0 /anc:1 /w:[ 1 1 1 ]
  and g32 (.I0(w29), .I1(w28), .Z(w30));   //: @(746,238) /sn:0 /w:[ 1 5 0 ]
  //: joint g27 (w24) @(529, 365) /w:[ 1 2 4 -1 ]
  buf g19 (.I(w20), .Z(w19));   //: @(600,437) /sn:0 /anc:1 /w:[ 1 0 ]
  and g38 (.I0(w35), .I1(w36), .Z(w33));   //: @(661,363) /sn:0 /w:[ 1 1 5 ]
  //: comment g6 /dolink:0 /link:"" @(22,11) /sn:0 /anc:1
  //: /line:"Dieses Tutorium f�hrt in spezielle Editiervorg�nge auf Leitungen ein."
  //: /end
  //: comment g53 /dolink:0 /link:"" @(726,534) /sn:0
  //: /line:"<---"
  //: /end
  //: comment g7 /dolink:0 /link:"" @(508,162) /sn:0 /anc:1
  //: /line:"<---"
  //: /end
  //: comment g9 /dolink:0 /link:"" @(26,30) /anc:1
  //: /line:"1) In TkGate ist ein besonderes \"Schwerkraftfeld\" "
  //: /line:"eingebaut. Kurze Leitungssegmente werden automatisch"
  //: /line:"bereinigt. Klicke auf den Draht am durch den Pfeil "
  //: /line:"gekennzeichneten Punkt in Bild 1 und bewege ihn, bis"
  //: /line:"er zu dem anderen vertikalen Leitungsabschnitt fast"
  //: /line:"ausgerichtet ist. Beim Ausl�ssen der Maustaste rasten"
  //: /line:"die beiden Segmente perfekt ausgerichtet ein."
  //: /line:""
  //: /line:"2) Tkgate l�scht automatisch Leitungsabschnitte, die "
  //: /line:"Schleifen bilden. Zur Demonstration w�hle das Ende der"
  //: /line:"Ausgangsleitung des XOR-Gatters in Bild 2 mit der linken"
  //: /line:"Maustaste aus. Ziehe das Ende nach oben direkt zum "
  //: /line:"Ausgang des Gatters und l�se die Maustaste aus. Diese"
  //: /line:"Automatik kann ausgeschaltet werden: Dr�cke beim "
  //: /line:"Bewegen von Dr�hten die \"ALT\"-Taste."
  //: /line:""
  //: /line:"3) TkGate ist auch in der Lage, unbenutzte "
  //: /line:"Verbindungspunkte automatisch zu l�schen. W�hle die"
  //: /line:"Kneifzange aus und schneide den Draht an der in Bild"
  //: /line:"3a angegebenen Stelle auf. Beachte, dass der L�tpunkt"
  //: /line:"automatisch entfernt wird. Ein Schnitt auf das freie"
  //: /line:"Ende in Bild 3b beseitigt dieses r�ckstandsfrei."
  //: /line:""
  //: /line:"4) Schalte zur�ck auf Bewegen/Verbinden und w�hle den "
  //: /line:"Eingang des untersten Puffers in Bild 4a aus, so da�"
  //: /line:"der L�tkolben erscheint. Bewege den Endpunkt in die"
  //: /line:"N�he der L�tstelle und l�se die Maustaste aus. Der"
  //: /line:"Draht wird mit der L�tstelle verbunden. Wiederhole die"
  //: /line:"Aktion in Bild 4b und l�se die Maustaste zwischen dem "
  //: /line:"AND-Gatter und der L�tstelle aus. Diesesmal wird eine"
  //: /line:"neue L�tstelle erzeugt."
  //: /line:""
  //: /line:"5) F�ge zum Ausgang des AND-Gatters in Bild 5 ein neues"
  //: /line:"Segment hinzu, um es mit dem gemeinsamen Eingang der"
  //: /line:"beiden Puffer zu verbinden. Klicke dazu mit der rechten"
  //: /line:"Maustaste auf das durch den Pfeil gekennzeichnete "
  //: /line:"Leitungssegment. W�hle dann \"Leitungssegment hinzuf�gen\""
  //: /line:"aus dem eingeblendeten Menu. Jetzt kann das Ende des"
  //: /line:"erzeugten Segments irgendwo mit dem Draht am Eingang"
  //: /line:"der beiden Puffer verbunden werden."
  //: /line:""
  //: /line:"6) W�hle die Leitung an den in den Bildern 6a und 6b"
  //: /line:"gekennzeichneten Punkten aus und ziehe sie nach links"
  //: /line:"hinter den Ausgangs-Punkt des AND-Gatters bzw. hinter"
  //: /line:"die Position des Verbindungspunktes. Im Fall des "
  //: /line:"AND-Gatters werden Segmente hinzugef�gt, damit der"
  //: /line:"die Leitung den Ausgang mit Sicherheit nach rechts "
  //: /line:"verl��t. Im Fall des L�tpunktes wird die"
  //: /line:"Position des Drahtes rund um diesen Verbindungspunkt"
  //: /line:"neu justiert. "
  //: /end
  //: joint g31 (w28) @(705, 286) /w:[ 2 4 1 -1 ]
  //: comment g20 /dolink:1 /link:"@T/create_tut.v" @(630,55) /sn:0 /anc:1
  //: /line:"Erzeugen einer Schaltung"
  //: /end
  //: frame g15 @(600,25) /sn:0 /anc:1 /wi:213 /ht:149 /tx:"Tutorien"
  and g39 (.I0(w13), .I1(w41), .Z(w42));   //: @(520,549) /sn:0 /anc:1 /w:[ 1 1 0 ]
  buf g48 (.I(w46), .Z(w47));   //: @(743,572) /sn:0 /w:[ 0 0 ]
  //: frame g43 @(624,224) /sn:0 /anc:1 /wi:160 /ht:85 /tx:"Bild 3b"
  buf g29 (.I(w23), .Z(w27));   //: @(560,393) /sn:0 /w:[ 1 0 ]
  and g25 (.I0(w10), .I1(w22), .Z(w24));   //: @(479,365) /sn:0 /w:[ 1 1 5 ]
  //: comment g17 /dolink:1 /link:"@T/sim_tut.v" @(630,130) /sn:0 /anc:1
  //: /line:"Schaltnetzsimulation"
  //: /end
  //: frame g52 @(612,509) /sn:0 /anc:1 /wi:189 /ht:73 /tx:"Bild 6b"
  //: frame g42 @(448,226) /sn:0 /anc:1 /wi:163 /ht:83 /tx:"Bild 3a"
  and g5 (.I0(w7), .I1(w9), .Z(w17));   //: @(497,438) /sn:0 /w:[ 1 1 1 ]
  //: comment g14 /dolink:1 /link:"@T/seqsim_tut.v" @(630,145) /sn:0 /anc:1
  //: /line:"Schaltwerkssimulation"
  //: /end
  and g47 (.I0(w43), .I1(w44), .Z(w46));   //: @(649,561) /sn:0 /w:[ 1 1 5 ]
  buf g44 (.I(w37), .Z(w38));   //: @(745,394) /sn:0 /w:[ 1 0 ]
  buf g36 (.I(w33), .Z(w34));   //: @(742,363) /sn:0 /w:[ 0 0 ]
  //: comment g24 /dolink:0 /link:"" @(491,449) /sn:0
  //: /line:"--->"
  //: /end
  //: comment g21 /dolink:1 /link:"@T/edit2_tut.v" @(630,85) /sn:0 /anc:1
  //: /line:"Editieren von Gruppen"
  //: /end
  //: frame g41 @(447,128) /sn:0 /anc:1 /wi:142 /ht:86 /tx:"Bild 2"
  buf g23 (.I(w20), .Z(w21));   //: @(600,475) /sn:0 /anc:1 /w:[ 0 0 ]
  //: comment g54 /dolink:0 /link:"" @(556,521) /sn:0 /anc:1
  //: /line:"<---"
  //: /end
  //: frame g40 @(442,34) /sn:0 /anc:1 /wi:147 /ht:86 /tx:"Bild 1"
  //: frame g46 @(449,419) /sn:0 /anc:1 /wi:190 /ht:75 /tx:"Bild 5"
  buf g45 (.I(w33), .Z(w39));   //: @(743,331) /sn:0 /w:[ 3 0 ]
  //: frame g35 @(627,319) /sn:0 /anc:1 /wi:159 /ht:88 /tx:"Bild 4b"
  buf g26 (.I(w24), .Z(w25));   //: @(561,334) /sn:0 /w:[ 3 0 ]
  //: comment g22 /dolink:0 /link:"" @(605,100) /sn:0 /anc:1
  //: /line:"->"
  //: /end
  and g0 (.I0(w1), .I1(w2), .Z(w3));   //: @(479,288) /sn:0 /w:[ 1 1 0 ]
  //: comment g12 /dolink:0 /link:"" @(552,63) /sn:0 /anc:1
  //: /line:"<---"
  //: /end
  //: comment g18 /dolink:1 /link:"@T/welcome_tut.v" @(630,40) /sn:0 /anc:1
  //: /line:"TkGate Einf�hrung"
  //: /end
  and g33 (.I0(w31), .I1(w32), .Z(w28));   //: @(652,286) /sn:0 /w:[ 1 1 0 ]
  //: comment g30 /dolink:0 /link:"" @(730,252) /sn:0 /anc:1
  //: /line:"|"
  //: /line:"v"
  //: /end
  buf g49 (.I(w46), .Z(w48));   //: @(741,523) /sn:0 /anc:1 /w:[ 3 0 ]

endmodule
