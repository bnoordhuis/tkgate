//: version "2.0"
//: property prefix = "_GG"
//: property title = "label.v"

//: /netlistBegin main
module main;    //: root_module
wire w6;    //: /sn:0 {0}(587,324)(587,339){1}
wire w7;    //: /sn:0 {0}(374,112)(389,112){1}
wire w4;    //: /sn:0 {0}(409,529)(424,529){1}
wire w0;    //: /sn:0 {0}(140,135)(155,135){1}
wire w3;    //: /sn:0 {0}(567,324)(567,339){1}
wire w1;    //: /sn:0 {0}(140,140)(155,140){1}
wire w8;    //: /sn:0 {0}(539,355)(554,355){1}
wire w2;    //: /sn:0 {0}(338,109)(353,109){1}
wire w11;    //: /sn:0 {0}(478,440)(478,455){1}
wire w12;    //: /sn:0 {0}(430,471)(445,471){1}
wire w10;    //: /sn:0 {0}(458,440)(458,455){1}
wire w13;    //: /sn:0 {0}(468,484)(468,499){1}
wire w5;    //: /sn:0 {0}(445,527)(460,527){1}
wire w9;    //: /sn:0 {0}(577,368)(577,383){1}
wire FOOBAR;    //: {0}(424,524)(-50:293,524)(293,384)(80:187,384)(187,304){1}
//: {2}(189,302)(234,302)(234,114)(353,114){3}
//: {4}(185,302)(175,302)(175,153)(186,153)(186,138)(176,138){5}
//: enddecls

  _GGMUX2 #(4, 2) g4 (.I0(w3), .I1(w6), .S(w8), .Z(w9));   //: @(577,355) /sn:0 /delay:" 4 2" /w:[ 1 1 1 0 ] /ss:0 /do:0
  //: joint g3 (FOOBAR) @(187, 302) /w:[ 2 -1 4 1 ]
  _GGAND2 #(3) g2 (.I0(w2), .I1(FOOBAR), .Z(w7));   //: @(364,112) /sn:0 /delay:" 3" /w:[ 1 3 0 ]
  _GGAND2 #(6) g1 (.I0(FOOBAR), .I1(w4), .Z(w5));   //: @(435,527) /sn:0 /w:[ 0 1 0 ]
  foo #(.B(42)) g6 ();   //: @(307, 278) /sz:(40, 40) /sn:0 /p:[ ]
  _GGMUX2 #(8, 8) g5 (.I0(w10), .I1(w11), .S(w12), .Z(w13));   //: @(468,471) /sn:0 /w:[ 1 1 1 0 ] /ss:0 /do:0
  _GGAND2 #(6) g0 (.I0(w0), .I1(w1), .Z(FOOBAR));   //: @(166,138) /sn:0 /w:[ 1 1 5 ]

endmodule
//: /netlistEnd

//: /hdlBegin foo
//: interface  /sz:(40, 40) /bd:[ ]
//: enddecls
module foo #(.A(8), .B(99)) (X,Y,Z);

endmodule
//: /hdlEnd
