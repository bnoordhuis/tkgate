//: version "2.0-b6"
//: property encoding = "euc-jp"
//: property locale = "ja"
//: property prefix = "_GG"
//: property title = "Welcome to TkGate Page"
//: property discardChanges = 1

`timescale 1ns/1ns

//: /netlistBegin PAGE1
module PAGE1;    //: root_module
//: enddecls

  //: comment g1 @(433,291) /sn:0 /R:14
  //: /line:"<a href=\"welcome.v\">TkGate�Υᥤ��Υڡ�������롣</a>"
  //: /end
  //: comment g0 @(434,49) /sn:0 /anc:1
  //: /line:"<a href=\"welcome.v\"><img src=\"biggatelogo.gif\"></a>"
  //: /end
  //: comment g18 @(10,10) /sn:0 /anc:1
  //: /line:"<h1>���塼�ȥꥢ��ξϤΰ���ɽ:</h1>"
  //: /line:""
  //: /line:"<h3><a href=\"create.v\">1. ��ϩ�κ���</a></h3> - Get started by creating a simple circuit."
  //: /line:""
  //: /line:"<h3><a href=\"gates.v\">2. �����Ȥ��Խ�</a></h3> - The basics of editing gates."
  //: /line:""
  //: /line:"<h3><a href=\"wires.v\">3. �磻����Խ�</a></h3> - The basics of editing wires."
  //: /line:""
  //: /line:"<h3><a href=\"group.v\">4. ���롼���Խ��ε�ǽ</a></h3> - Operate on groups of gates."
  //: /line:""
  //: /line:"<h3><a href=\"modules.v\">5. �桼�����⥸�塼��</a></h3> - Using modules in your circuit."
  //: /line:""
  //: /line:"<h3><a href=\"advanced.v\">6. Advanced Editing Techniques</a></h3> - Learn advanced editing tricks."
  //: /line:""
  //: /line:"<h3><a href=\"combinational1.v\">7. �ȹ礻��ϩ�Υ��ߥ�졼�����</a></h3> - Simulate a circuit with"
  //: /line:"    combinational logic."
  //: /line:""
  //: /line:"<h3><a href=\"sequential1.v\">8. �����ϩ�Υ��ߥ�졼�����</a></h3> - Simulate a circuit with"
  //: /line:"    sequential logic."
  //: /line:""
  //: /line:"<h3><a href=\"verilog.v\">9. �ƥ�����Verilog</a></h3> - Create modules with textual Verilog descriptions."
  //: /line:""
  //: /line:"<h3><a href=\"options.v\">10. TkGate�Υ��ץ����</a></h3> - Customize TkGate to suit your tastes."
  //: /line:""
  //: /line:""
  //: /line:""
  //: /end

endmodule
//: /netlistEnd


`timescale 1ns/1ns

