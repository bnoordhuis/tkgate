//: version "2.0"
//: property title = "create_tut.v"
//: property useExtBars = 0
//: property discardChanges = 1

module main;    //: root_module
wire w6;    //: /sn:0 {0}(232,502)(177,502){1}
//: {2}(175,500)(175,466)(187,466){3}
//: {4}(173,502)(141,502){5}
wire w7;    //: /sn:0 {0}(253,500)(263,500){1}
wire w2;    //: /sn:0 {0}(187,461)(141,461){1}
wire w5;    //: /sn:0 {0}(232,497)(218,497)(218,464)(208,464){1}
//: enddecls

  or g4 (.I0(w5), .I1(w6), .Z(w7));   //: @(243,500) /sn:0 /anc:1 /w:[ 0 0 0 ]
  //: comment g8 @(248,476) /anc:1
  //: /line:"OR������"
  //: /end
  //: comment g61 @(622,100) /sn:0
  //: /line:"<a href=\"@T/edwire_tut.v\">�磻����Խ�</a>"
  //: /end
  //: frame g13 @(412,372) /sn:0 /wi:381 /ht:177 /tx:"��ϩ�򤳤���˺������Ʋ�����"
  and g3 (.I0(w2), .I1(w6), .Z(w5));   //: @(198,464) /sn:0 /anc:1 /w:[ 0 3 1 ]
  //: switch g2 (w6) @(124,502) /sn:0 /anc:1 /w:[ 5 ] /st:0
  //: switch g1 (w2) @(124,461) /sn:0 /anc:1 /w:[ 1 ] /st:0
  //: comment g16 @(622,115) /sn:0
  //: /line:"<a href=\"@T/module_tut.v\">�⥸�塼��λȤ���</a>"
  //: /end
  //: comment g10 @(11,205) /anc:1
  //: /line:"5) AND�����Ȥ�OR�����Ȥ�Ʊ���ͤ���ĤΥ����å���������Ʋ��������κ����ϥ�˥塼�Ρ�I/O��"
  //: /line:"���֥�˥塼�ΡΥ����å��Ϥ�����ǡ����ϡ������ܡ��ɡ����硼�ȥ��åȤ�\"s\"�򲡤��Ʋ�������"
  //: /line:""
  //: /line:"6) ���ƥå�4�򷫤��֤��ơ���Υ����å��ν��Ϥ�AND�����Ȥξ�ν��Ϥ���³���Ʋ�������"
  //: /line:""
  //: /line:"7) ���ƥå�4�򷫤��֤��ơ����Υ����å��ν��Ϥ�OR�����Ȥβ��ν��Ϥ���³���Ʋ�������"
  //: /line:""
  //: /line:"8) AND�����Ȥβ������Ϥ򥯥�å����ơ��Ϥ�����Ƥ�Ф������Υ����å���OR�����Ȥδ֤�"
  //: /line:"�磻��ο���˥ɥ�å����ơ��ޥ����ܥ����Υ���Ʋ���������³������������ޤ���"
  //: /end
  //: comment g6 @(101,427) /anc:1
  //: /line:"�����å�"
  //: /end
  //: comment g7 @(192,436) /anc:1
  //: /line:"AND������"
  //: /end
  //: comment g9 @(12,9) /anc:1
  //: /line:"1) ���Υ��塼�ȥꥢ��Ǥϡ����˼����Ƥ���Τ�Ʊ���ͤʲ�ϩ��������롣������"
  //: /line:"����Ȣ����˺������Ʋ��������ޤ����ޥ����α��ܥ����AND�����Ȥΰ��֤������"
  //: /line:"������������å��������֤�X���ȡκ����ϥ�˥塼������ޤ���"
  //: /line:""
  //: /line:"2) ���줫�顢�κ����ϥ�˥塼�ΡΥ����ȡϥ��֥�˥塼�Ρ�AND�Ϥ�����ǲ�������"
  //: /line:"��˥塼���С������ϥ����ܡ��ɡ����硼�ȥ��åȤ�\"a\"��Ȥ��ޤ���"
  //: /line:""
  //: /line:"3) ���ƥå�1��2�򷫤��֤���, OR�����Ȥ�AND�����Ȥα����ΰ��֤˺������Ʋ�������"
  //: /line:"��˥塼���С������ϥ����ܡ��ɥ��硼�ȡ����åȤ�\"o\"��Ȥ��ޤ���"
  //: /line:""
  //: /line:"4) AND�����Ȥν��ϤΥ磻�����ü��ޥ����κ��ܥ���ǥ���å����ơ��ܥ���򲡤�"
  //: /line:"���ޤޤˤ��ޤ����ޥ������������뤬�Ϥ�����Ƥ��Ѥ��ޤ����磻���OR�����Ȥ�"
  //: /line:"������Ϥޤǥɥ�å����ƥޥ������ܥ����Υ���ȡ��磻�䤬��³����ޤ���"
  //: /end
  //: frame g15 @(600,25) /sn:0 /wi:224 /ht:149 /tx:"���塼�ȥꥢ��"
  //: comment g20 @(622,55) /sn:0 /anc:1
  //: /line:"��ϩ�κ���"
  //: /end
  //: comment g17 @(622,130) /sn:0
  //: /line:"<a href=\"@T/sim_tut.v\">�ȹ礻��ϩ�Υ��ߥ�졼�����</a>"
  //: /end
  //: joint g5 (w6) @(175, 502) /anc:1 /w:[ 1 2 4 -1 ]
  //: comment g14 @(622,145) /sn:0
  //: /line:"<a href=\"@T/seqsim_tut.v\">�����ϩ�Υ��ߥ�졼�����</a>"
  //: /end
  //: comment g21 @(622,85) /sn:0
  //: /line:"<a href=\"@T/edit2_tut.v\">���롼�פ��Խ���ǽ</a>"
  //: /end
  //: comment g0 @(622,70) /sn:0
  //: /line:"<a href=\"@T/edit1_tut.v\">���ܤ��Խ��⡼��</a>"
  //: /end
  //: comment g22 @(605,55) /sn:0
  //: /line:"->"
  //: /end
  //: comment g18 @(622,40) /sn:0
  //: /line:"<a href=\"@T/welcome_tut.v\">TkGate�ξҲ�</a>"
  //: /end

endmodule
