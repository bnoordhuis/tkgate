//: version "2.0"
//: property title = "edit2_tut.v"
//: property useExtBars = 0
//: property discardChanges = 1

module main;    //: root_module
wire w3;    //: /sn:0 {0}(756,264)(679,264){1}
wire w1;    //: /sn:0 {0}(756,259)(712,259)(712,224)(679,224){1}
wire w2;    //: /sn:0 {0}(679,302)(689,302){1}
wire w5;    //: /sn:0 {0}(777,262)(787,262){1}
//: enddecls

  and g4 (.I0(w1), .I1(w3), .Z(w5));   //: @(767,262) /sn:0 /w:[ 0 0 0 ]
  //: comment g61 /dolink:1 /link:"@T/edwire_tut.v" @(622,100) /sn:0
  //: /line:"�磻����Խ�"
  //: /end
  //: switch g3 (w2) @(662,302) /sn:0 /w:[ 0 ] /st:0
  //: switch g2 (w3) @(662,264) /sn:0 /w:[ 1 ] /st:0
  //: switch g1 (w1) @(662,224) /sn:0 /w:[ 1 ] /st:0
  //: frame g11 @(434,347) /sn:0 /anc:1 /wi:373 /ht:230 /tx:"�����Ȥ򤳤���˥��ԡ�����"
  //: comment g16 /dolink:1 /link:"@T/module_tut.v" @(622,115) /sn:0
  //: /line:"�⥸�塼��λȤ���"
  //: /end
  //: frame g10 @(22,347) /sn:0 /anc:1 /wi:394 /ht:227 /tx:"�����Ȥ򤳤���˰�ư����"
  //: comment g6 /dolink:1 /link:"@T/edit1_tut.v" @(622,70) /sn:0
  //: /line:"���ܤ��Խ��⡼��"
  //: /end
  //: comment g9 /dolink:0 /link:"" @(607,452) /sn:0
  //: /line:""
  //: /end
  //: comment g7 /dolink:0 /link:"" @(634,193) /sn:0
  //: /line:""
  //: /end
  //: frame g15 @(600,25) /sn:0 /wi:224 /ht:149 /tx:"���塼�ȥꥢ��"
  //: comment g20 /dolink:1 /link:"@T/create_tut.v" @(622,55) /sn:0
  //: /line:"��ϩ�κ���"
  //: /end
  //: comment g17 /dolink:1 /link:"@T/sim_tut.v" @(622,130) /sn:0
  //: /line:"�ȹ礻��ϩ�Υ��ߥ�졼�����"
  //: /end
  //: comment g5 /dolink:0 /link:"" @(38,36) /anc:1
  //: /line:"1) �ޥ������ܥ���Ǳ��ˤ����ϩ�κ���򥯥�å����ơ�Ȣ����ϩ������"
  //: /line:"�ޤ�ޤǥޥ����򱦲��إɥ�å����ơ��ܥ����Υ���Ʋ�������"
  //: /line:"�����Ȥ����򤵤졢������ɽ������ޤ������򤵤�Ƥ��륲���Ȥν����"
  //: /line:"���쥯�����Ȥ����ޤ���"
  //: /line:""
  //: /line:"2) �����ȤΤɤ줫�򥯥�å����ơ֥����Ȥ򤳤���˰�ư����פȽ񤤤Ƥ���"
  //: /line:"������Ȣ����˰�ư���ƤߤƲ������������Ȥ�磻��Τʤ���򥯥�å������"
  //: /line:"���쥯�����ϲ������ޤ���"
  //: /line:""
  //: /line:"3) AND�����Ȥ����򤷤ơ��ޥ������ܥ���򲡤��������Ϥ��ɲáפ����򤷤�"
  //: /line:"�����������줫��AND�����Ȥ��ɲä��줿�磻��򲼤Υ����å�����³���Ʋ�������"
  //: /line:""
  //: /line:"4) ���ƥå�1�˽񤤤Ƥ����ͤ����ƤΥ����Ȥ����򤷤Ƥ����Ʋ����������줫��"
  //: /line:"���Խ��ץ�˥塼�Ρ֥��ԡ��פ����򤷡��ޥ������ܥ���ǡ֥����Ȥ򤳤����"
  //: /line:"���ԡ�����פȽ񤤤Ƥ���������Ȣ�ο���򥯥�å����ơ����Խ��ץ�˥塼��"
  //: /line:"��ĥ���դ��פ����򤷤Ʋ������������ȤΥ��쥯����󤬥��ԡ�����ޤ������쥯"
  //: /line:"����󤬤�������ǥ꡼�ȡ������򲡤��ȡ����쥯�����Υ����Ȥ��������ޤ���"
  //: /line:""
  //: /line:"5) ����ȥ��롦�����򲡤��ʤ��顢�����Ȥ򥯥�å�����ȡ������Ȥ��Ĥ���"
  //: /line:"���쥯�������ɲä��뤳�Ȥ�����ޤ���"
  //: /end
  //: comment g14 /dolink:1 /link:"@T/seqsim_tut.v" @(622,145) /sn:0
  //: /line:"�����ϩ�Υ��ߥ�졼�����"
  //: /end
  //: comment g21 /dolink:0 /link:"@T/edit2_tut.v" @(622,85) /sn:0 /anc:1
  //: /line:"���롼�פ��Խ���ǽ"
  //: /end
  //: comment g0 /dolink:0 /link:"" @(26,17) /anc:1
  //: /line:"���Υ��塼�ȥꥢ��ϥ��롼���Խ��ε�ǽ��Ҳ𤹤롣"
  //: /end
  //: comment g22 /dolink:0 /link:"" @(605,85) /sn:0
  //: /line:"->"
  //: /end
  //: comment g18 /dolink:1 /link:"@T/welcome_tut.v" @(622,40) /sn:0
  //: /line:"TkGate�ξҲ�"
  //: /end

endmodule
