//: version "2.0"
//: property title = "notes.v"

module main;    //: root_module
//: enddecls

  //: comment g1 /dolink:1 /link:"@T/welcome_tut.v" @(611,27) /sn:0
  //: /line:"Return to welcome."
  //: /end
  //: comment g0 /dolink:0 /link:"" @(42,57) /sn:0
  //: /line:"* Make sure interface in library matches interfaces used in circuit."
  //: /line:"* Add HDL module type."
  //: /line:"* HTML tags in comments instead of all-or-nothing hyperlink."
  //: /line:"* How about a simulator selection dialog box with options for switches to include, etc."
  //: /line:"* Bitmap symbol editor for libraries"
  //: /line:"* HDL modules"
  //: /line:"* Current module's interface shown in lower left box."
  //: /line:""
  //: /line:"BUGS:"
  //: /line:"* Landscape printing with A4 paper."
  //: /line:"* Lack of editing on edit interfaces screen."
  //: /line:"* Mysterious double modules on interface screen in welcome_tut.v"
  //: /line:"* Ctl-D duplicate a gate, then double click.  prop box doesn't open."
  //: /line:""
  //: /line:"TO DO:"
  //: /line:""
  //: /line:"* Finish module interface generator"
  //: /line:"* Convert port box to use SpreadSheet"
  //: /line:"* Verilog Modules"
  //: /line:"* Custom Module Symbols"
  //: /line:"* Dialog box images"
  //: /line:"* Japanese messages.ja"
  //: /line:""
  //: /end

endmodule
